LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY ram8 IS
    PORT (
        input : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        address : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        load : IN STD_LOGIC;
        clk : IN STD_LOGIC;
        output : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
    );
END ENTITY ram8;

ARCHITECTURE ram8_arch OF ram8 IS
    -- load signals for each register
    SIGNAL load_0 : STD_LOGIC;
    SIGNAL load_1 : STD_LOGIC;
    SIGNAL load_2 : STD_LOGIC;
    SIGNAL load_3 : STD_LOGIC;
    SIGNAL load_4 : STD_LOGIC;
    SIGNAL load_5 : STD_LOGIC;
    SIGNAL load_6 : STD_LOGIC;
    SIGNAL load_7 : STD_LOGIC;
    -- output signals for each register
    SIGNAL output_0 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL output_1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL output_2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL output_3 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL output_4 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL output_5 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL output_6 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL output_7 : STD_LOGIC_VECTOR(15 DOWNTO 0);
BEGIN
    -- dmux for load signals
    load_decoder : ENTITY work.decoder8way(decoder8way_arch)
        PORT MAP(
            sel => address,
            out_0 => load_0,
            out_1 => load_1,
            out_2 => load_2,
            out_3 => load_3,
            out_4 => load_4,
            out_5 => load_5,
            out_6 => load_6,
            out_7 => load_7
        );

    -- getting the outputs from the registers
    register_0 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_0, clk => clk, output => output_0);
    register_1 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_1, clk => clk, output => output_1);
    register_2 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_2, clk => clk, output => output_2);
    register_3 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_3, clk => clk, output => output_3);
    register_4 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_4, clk => clk, output => output_4);
    register_5 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_5, clk => clk, output => output_5);
    register_6 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_6, clk => clk, output => output_6);
    register_7 : ENTITY work.regist(regist_arch)
        PORT MAP (input => input, load => load_7, clk => clk, output => output_7);

    -- selecting the output
    mux8way16_comp : ENTITY work.mux8way16(mux8way16_arch)
        PORT MAP(
            a => output_0,
            b => output_1,
            c => output_2,
            d => output_3,
            e => output_4,
            f => output_5,
            g => output_6,
            h => output_7,
            sel => address,
            output => output
        );

END ARCHITECTURE ram8_arch;